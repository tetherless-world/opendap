// This CDL file is a mockup for how to represent the following tabular LiDAR data:
//
// lat lon alt intensity category(Ground=2;Low-Vegitation=3;Unclassified=1;Water=9)
// 414783.24 3741669.72 40.32 26 Water
// 414782.09 3741669.31 40.44 3 Water
// 414782.73 3741670.04 40.40 10 Water
// 414782.03 3741670.63 40.28 26 Water
// 414781.51 3741671.03 40.34 22 Water
//
// NOTE: We're assuming that the non-uniform lat/long becomes uniformly gridded.
//       This doesn't make much sense for LiDAR data.
//
//3> <> prov:specializationOf 
//3>   <https://github.com/tetherless-world/opendap/blob/master/data/source/usgs-gov/earthexplorer/version/disneyland-2014-Jan-31/manual/CA_OrangeCo_2011_000402.sample.cdl>;
//3>    prov:wasDerivedFrom <http://www.unidata.ucar.edu/software/netcdf/workshops/2010/apis_examples/ExampleDataset2D.html>;
//3> .

netcdf disneyland_lidar {

dimensions:
   latitude  = 5 ;
   longitude = 1 ;

variables:
   float latitude(latitude) ;
      latitude:units = "?" ;
   float longitude(longitude) ;
      longitude:units = "?" ;
   float altitude(latitude, longitude) ;
      altitude:units = "?" ;
   float intensity(latitude, longitude) ;
      intensity:units = "?" ;
   int category(latitude, longitude) ;

data:
   // This sets up the grid that we don't actually want to assume.
   // ERROR: We're rounding to get to a grid.
   latitude  = 414781.5, 414782, 414782.5, 414783, 414783.5 ; 
   // ERROR: We're squashing to get to a grid.
   longitude = 3741670 ; 

   altitude =
      40.32,
      40.44,
      40.40,
      40.28,
      40.34 ;

   intensity =
      26,
      3,
      10,
      26,
      22 ;

   category =
      9,
      9,
      9,
      9,
      9 ;
}
