// This CDL file is a mockup for how to represent the following tabular data:
//
// lat lon alt intensity category;Ground=2 Low Vegitation=3 Unclassified=1 Water=9
// 414783.24 3741669.72 40.32 26 Water
// 414782.09 3741669.31 40.44 3 Water
// 414782.73 3741670.04 40.40 10 Water
// 414782.03 3741670.63 40.28 26 Water
// 414781.51 3741671.03 40.34 22 Water
//
// NOTE: We're assuming that the non-uniform lat/long becomes uniformly gridded.
//       This doesn't make much sense for LiDAR data.
//
//3> <> prov:specializationOf 
//3>   <https://github.com/tetherless-world/opendap/blob/master/data/source/usgs-gov/earthexplorer/version/disneyland-2014-Jan-31/manual/CA_OrangeCo_2011_000402.sample.cdl>;
//3>    prov:wasDerivedFrom <http://www.unidata.ucar.edu/software/netcdf/workshops/2010/apis_examples/ExampleDataset2D.html>;
//3> .

netcdf disneyland_lidar {

dimensions:
   latitude  = 6 ;
   longitude = 12 ;

variables:
   float latitude(latitude) ;
      latitude:units = "?" ;
   float longitude(longitude) ;
      longitude:units = "?" ;
   float altitude(latitude, longitude) ;
      altitude:units = "?" ;
   float intensity(latitude, longitude) ;
      intensity:units = "?" ;

data:
   // This sets up the grid that we don't actually want to assume.
   latitude  = 25, 30, 35, 40, 45, 50 ;
   longitude = -125, -120, -115, -110, -105, -100, -95, -90, -85, -80, -75, -70 ;

   altitude =
      900, 906, 912, 918, 924, 930, 936, 942, 948, 954, 960, 966,
      901, 907, 913, 919, 925, 931, 937, 943, 949, 955, 961, 967,
      902, 908, 914, 920, 926, 932, 938, 944, 950, 956, 962, 968,
      903, 909, 915, 921, 927, 933, 939, 945, 951, 957, 963, 969,
      904, 910, 916, 922, 928, 934, 940, 946, 952, 958, 964, 970,
      905, 911, 917, 923, 929, 935, 941, 947, 953, 959, 965, 971 ;

   intensity =
      9, 10.5, 12, 13.5, 15, 16.5, 18, 19.5, 21, 22.5, 24, 25.5,
      9.25, 10.75, 12.25, 13.75, 15.25, 16.75, 18.25, 19.75, 21.25, 22.75, 24.25, 25.75,
      9.5, 11, 12.5, 14, 15.5, 17, 18.5, 20, 21.5, 23, 24.5, 26,
      9.75, 11.25, 12.75, 14.25, 15.75, 17.25, 18.75, 20.25, 21.75, 23.25, 24.75, 26.25,
      10, 11.5, 13, 14.5, 16, 17.5, 19, 20.5, 22, 23.5, 25, 26.5,
      10.25, 11.75, 13.25, 14.75, 16.25, 17.75, 19.25, 20.75, 22.25, 23.75, 25.25, 26.75 ;
}
